module top(input clk,
	input  dout,			
	output adc_cs_n,			
	output din,					
	output adc_sck,
	output [3:0]dc,
	output l_w,
	output r_w,
	output c_w,
	output tx,
	output [8:0] rgb_w,
	input freq_color,
	output s2,
	output s3,
	output reg [1:0]turn_w
	);
	
reg [32:0] ct_pwm = 0;
wire l;
wire r;
wire c;
reg [2:0] rgb_w1[3];
reg [3:0]dc_r ='b0000;
//////////////////////////////////////////////
adc_control(.clk_50(clk),
					.dout(dout),
					.adc_cs_n(adc_cs_n),
					.din(din),
					.adc_sck(adc_sck),
					.l(l),
					.r(r),
					.c(c));

//////////////////////////////////////////////

////////////////////////////////////////////////
wire[2:0] rgb;
top_color(.clk(clk),
				.s2(s2),
				.s3(s3),
				.ip_signal(freq_color),
				.color(rgb));


///////////////////////////////////////////////

//uart
////////////////////////////////////////////	
integer msg_index=0;
reg transmit =0;
reg [1:0] node_t = 'b01;
wire uart_done;
reg [64:0] str[3];
integer msg_jndex =0;
reg [63:0]tstr;
uart(.clk(clk),
		.transmit(transmit),
		.str(tstr),
		.tx(tx),
		.done(uart_done));
		
//uart initial//		
initial
begin
str[0]="GBI3-D-#";
str[1]="GBI2-W-#";
str[2]="GBI1-M-#";
end	



////////////////////////////////////////////////
	

//////////////////////////////////////////////
reg p_start=0;
reg [4:0]s_node;
reg [4:0]e_node;
wire p_done;
wire [10*2-1:0] final_path;
path_planner(.clk(clk),
				 .start(p_start),
				 .s_node(s_node),
				 .e_node(e_node),
				 .done(p_done),
				 .final_path(final_path));
				 
				 
initial
begin
s_node = 0;
e_node = 3;
end
////////////////////////////////////////////
	
integer ct =0;
integer state=1;
reg [19:0] temp_path;
reg [32:0]delay = 0;
integer i =0;
integer nn = 0;
integer next_node[2];
integer line_follow_state; 
integer turn =0;
integer st = 1;
reg [1:0]ledi=0;
reg end_of_run = 0;
////////////////////////////////////////////
	
initial
begin
next_node[0]=8;
next_node[1]=14;
end
always @(posedge clk)
begin
if(transmit ==1)
transmit=0;
case(st)
5:
begin
dc_r = 4'b0;
case(state)
1:
begin
if(ct<100)
p_start=1;
else
begin
ct=0;
p_start =0;
state=2;
end
ct = ct+1;
end
2:
begin
if(p_done ==1)
begin
temp_path <= final_path;
state = 3;
end
end
3:
begin
delay = delay +1;
if(delay == 'd50000000)
begin
delay = 0;
turn_w[0] = temp_path[i];
turn_w[1] = temp_path[i+1];
i=i+2;
if(turn_w[0]==1 && turn_w[1]==0)
turn = 6;
if(turn_w[0]==0 && turn_w[1]==1)
turn =7;
if(turn_w[0]==1 && turn_w[1]==1)
turn =8;
if(turn_w[0] ==0 && turn_w[1]==0)
begin
st=4;
turn = 4;
if(e_node ==14)
begin
end_of_run =1;
st =4;                  ////////////////end of run//////////////////
state = 4;
end
else
begin
i=0;
state =1;
s_node = e_node;
e_node = next_node[nn];
nn = nn+1;
end
end
if(st !=4)
st = 3;
end
end
endcase
end


3:
begin
case(turn)
0:
dc_r[3:0]=4'b0;

4:											//u-turn
begin

dc_r[1:0] = 'b10;
dc_r[3:2] = 'b10;


end
5:											//back
begin
dc_r[1:0] = 'b01;
dc_r[3:2] = 'b10;
end
6:
begin
dc_r[1:0] = 'b00;
dc_r[3:2] = 'b01;
end
7:
begin
dc_r[1:0] = 'b10;
dc_r[3:2] = 'b00;
end


8:
begin
dc_r[1:0]='b10;
dc_r[3:2]='b01;
end
endcase
if(l==1 && c==0 && r==1)
begin
st = 1;        ///follow line
line_follow_state =1;
turn =0;       ///dead state of turn
end
end

4:
begin
rgb_w1[ledi] = rgb;
if(rgb_w1[ledi] == 'b001)
tstr = str[1];
if(rgb_w1[ledi] == 'b100)
tstr = str[2];
if(rgb_w1[ledi] == 'b010)
tstr = str[0];
ledi = ledi+'d1;
transmit = 1;
st=3;
if(end_of_run==1)
st=6;
end






1:                   ////////////////simple line following case///////////////////
begin
st = 1;
ct_pwm = ct_pwm +1;
if(ct_pwm=='d999999)ct_pwm=0;

if(l==0 && r==1)
begin
line_follow_state=2;
end

else if(l==1 && r==0)
begin
line_follow_state=3;
end
else if(l==1 && r==1 && c==0)
begin
line_follow_state =1;
end
else if(l==0 && r==0 && c==0)
begin
line_follow_state =0;
st =5;            ///on node go to delay line_follow_state.
end
 
if(ct_pwm<'d600000)
begin

case (line_follow_state)
0:											//stop
begin
dc_r[3:0] = 'b0;
end
1:                               //follow line
begin
dc_r[1:0] = 'b10;
dc_r[3:2] = 'b01;
end
2:                               //left turn
begin
dc_r[1:0] = 'b10;
dc_r[3:2] = 'b00;
end
3:											//right turn
begin
dc_r[1:0] = 'b00;
dc_r[3:2] = 'b01;
end

endcase
end
end                 ///////////////////line followning case ends here.../////////////






endcase
end
	
	
assign dc = dc_r;
assign l_w = l;
assign r_w = r;
assign c_w  =c;
assign rgb_w[2:0] = rgb_w1[0];
assign rgb_w[5:3] = rgb_w1[1];
assign rgb_w[8:6] = rgb_w1[2];

endmodule
